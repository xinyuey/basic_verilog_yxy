library verilog;
use verilog.vl_types.all;
entity spi_master_tb is
end spi_master_tb;
